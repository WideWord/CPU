
module SPICtl(
	input clk,
	input reset,
	
	output spi_clk,
	output spi_cmd,
	input spi_data,
	output spi_cs
	
);

endmodule
